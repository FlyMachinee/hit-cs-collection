module ram_top (
    input         clk,
    input  [15:0] ram_addr,
    input  [31:0] ram_wdata,
    input         ram_wen,
    output [31:0] ram_rdata
);

  block_ram block_ram (
      .clka (clk),
      .wea  (ram_wen),
      .addra(ram_addr),
      .dina (ram_wdata),
      .douta(ram_rdata)
  );
endmodule
